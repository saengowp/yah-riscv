00007137
00007437
00003517
50c50513
00050067
fd010113
02812623
03010413
fca42e23
fcb42c23
0a40006f
00004797
80478793
0007a783
0007c783
fef407a3
fef44783
0047d793
fef40723
fef44783
00f7f793
fef406a3
fed44783
00178793
0ff7f793
00f7f793
fef40623
fec44703
fee44783
00f71463
0540006f
00003797
7b478793
0007a703
fed44783
02078793
00f707b3
fdc42703
00074703
00e78023
00003797
79078793
0007a783
fec44703
00e78023
fdc42783
00178793
fcf42e23
fd842783
fff78793
fcf42c23
fd842783
f4079ee3
00000013
00000013
02c12403
03010113
00008067
fe010113
00812e23
02010413
00003797
73c78793
0007a783
0017c783
fef407a3
fef44783
00f7f793
fef407a3
fef44703
00003797
71c78793
0007a783
fcf708e3
00003797
70878793
0007a703
00003797
70078793
0007a783
01078793
00f707b3
0007c783
fef40723
00003797
6e478793
0007a783
00178793
00f7f713
00003797
6d078793
00e7a023
fee44783
00078513
01c12403
02010113
00008067
fd010113
02812623
03010413
fca42e23
fe042623
01c0006f
fec42783
00178793
fef42623
fdc42783
00178793
fcf42e23
fdc42783
0007c783
fe0790e3
fec42783
00078513
02c12403
03010113
00008067
fb010113
04812623
05010413
faa42e23
fe042623
0240006f
fec42783
00279793
ff078793
008787b3
fc07ae23
fec42783
00178793
fef42623
fec42703
00700793
fce7dce3
fbc42783
fcc42303
fd042883
fd442803
fd842503
fdc42583
fe042603
fe442683
fe842703
0067a023
0117a223
0107a423
00a7a623
00b7a823
00c7aa23
00d7ac23
00e7ae23
fbc42503
04c12403
05010113
00008067
fb010113
04112623
04812423
04912223
05212023
05010413
faa42e23
00058493
00060913
fcc40793
00078513
f3dff0ef
fe042623
0dc0006f
fec42783
00279793
00f487b3
0007a703
fec42783
00279793
00f907b3
0007a783
00f70733
fec42783
00279793
ff078793
008787b3
fdc7a783
00f70733
fec42783
00279793
ff078793
008787b3
fce7ae23
fec42783
00279793
ff078793
008787b3
fdc7a703
ffff07b7
00f777b3
06078063
fec42783
00279793
ff078793
008787b3
fdc7a703
ffff07b7
fff7c793
00f77733
fec42783
00279793
ff078793
008787b3
fce7ae23
fec42703
00700793
02f70063
fec42783
00178793
00279793
ff078793
008787b3
00100713
fce7ae23
fec42783
00178793
fef42623
fec42703
00700793
f2e7d0e3
fbc42783
fcc42303
fd042883
fd442803
fd842503
fdc42583
fe042603
fe442683
fe842703
0067a023
0117a223
0107a423
00a7a623
00b7a823
00c7aa23
00d7ac23
00e7ae23
fbc42503
04c12083
04812403
04412483
04012903
05010113
00008067
fb010113
04112623
04812423
04912223
05212023
05010413
faa42e23
00058493
00060913
fcc40793
00078513
dc1ff0ef
fe042623
0dc0006f
fec42783
00279793
00f487b3
0007a703
fec42783
00279793
00f907b3
0007a783
40f70733
fec42783
00279793
ff078793
008787b3
fdc7a783
40f70733
fec42783
00279793
ff078793
008787b3
fce7ae23
fec42783
00279793
ff078793
008787b3
fdc7a703
ffff07b7
00f777b3
06078063
fec42783
00279793
ff078793
008787b3
fdc7a703
ffff07b7
fff7c793
00f77733
fec42783
00279793
ff078793
008787b3
fce7ae23
fec42703
00700793
02f70063
fec42783
00178793
00279793
ff078793
008787b3
00100713
fce7ae23
fec42783
00178793
fef42623
fec42703
00700793
f2e7d0e3
fbc42783
fcc42303
fd042883
fd442803
fd842503
fdc42583
fe042603
fe442683
fe842703
0067a023
0117a223
0107a423
00a7a623
00b7a823
00c7aa23
00d7ac23
00e7ae23
fbc42503
04c12083
04812403
04412483
04012903
05010113
00008067
f5010113
0a112623
0a812423
0a912223
0b212023
0b010413
faa42e23
00058493
00060913
fcc40793
00078513
c45ff0ef
fe042623
1bc0006f
fec42783
41f7d713
00f77713
00f707b3
4047d793
00279793
00f907b3
0007a783
fec42703
00f77713
00100693
00e69733
00e7f7b3
0e078063
f9040313
fcc42883
fd042803
fd442503
fd842583
fdc42603
fe042683
fe442703
fe842783
f7142823
f7042a23
f6a42c23
f6b42e23
f8c42023
f8d42223
f8e42423
f8f42623
0004a883
0044a803
0084a503
00c4a583
0104a603
0144a683
0184a703
01c4a783
f5142823
f5042a23
f4a42c23
f4b42e23
f6c42023
f6d42223
f6e42423
f6f42623
f5040713
f7040793
00070613
00078593
00030513
c01ff0ef
f9042883
f9442803
f9842503
f9c42583
fa042603
fa442683
fa842703
fac42783
fd142623
fd042823
fca42a23
fcb42c23
fcc42e23
fed42023
fee42223
fef42423
0004a883
0044a803
0084a503
00c4a583
0104a603
0144a683
0184a703
01c4a783
f5142823
f5042a23
f4a42c23
f4b42e23
f6c42023
f6d42223
f6e42423
f6f42623
0004a883
0044a803
0084a503
00c4a583
0104a603
0144a683
0184a703
01c4a783
f7142823
f7042a23
f6a42c23
f6b42e23
f8c42023
f8d42223
f8e42423
f8f42623
f7040713
f5040793
00070613
00078593
00048513
b29ff0ef
fec42783
00178793
fef42623
fec42703
07f00793
e4e7d0e3
fbc42783
fcc42303
fd042883
fd442803
fd842503
fdc42583
fe042603
fe442683
fe842703
0067a023
0117a223
0107a423
00a7a623
00b7a823
00c7aa23
00d7ac23
00e7ae23
fbc42503
0ac12083
0a812403
0a412483
0a012903
0b010113
00008067
ff010113
00812623
00912423
01010413
00050493
01c4a783
00179713
ffff07b7
00f777b3
00078513
00c12403
00812483
01010113
00008067
fb010113
04812623
04912423
05010413
faa42e23
00058493
0004a883
0044a803
0084a503
00c4a583
0104a603
0144a683
0184a703
01c4a783
fd142623
fd042823
fca42a23
fcb42c23
fcc42e23
fed42023
fee42223
fef42423
fe042623
0ec0006f
fec42783
00279793
ff078793
008787b3
fdc7a783
0017d713
fec42783
00279793
ff078793
008787b3
fce7ae23
fec42703
00700793
04f70e63
fec42783
00279793
ff078793
008787b3
fdc7a703
fec42783
00178793
00279793
ff078793
008787b3
fdc7a783
00f79693
000107b7
fff78793
00f6f7b3
00f76733
fec42783
00279793
ff078793
008787b3
fce7ae23
0500006f
fec42783
00279793
ff078793
008787b3
fdc7a703
fec42783
00279793
ff078793
008787b3
fdc7a783
00179693
000087b7
00f6f7b3
00f76733
fec42783
00279793
ff078793
008787b3
fce7ae23
fec42783
00178793
fef42623
fec42703
00700793
f0e7d8e3
fbc42783
fcc42303
fd042883
fd442803
fd842503
fdc42583
fe042603
fe442683
fe842703
0067a023
0117a223
0107a423
00a7a623
00b7a823
00c7aa23
00d7ac23
00e7ae23
fbc42503
04c12403
04812483
05010113
00008067
ed010113
12112623
12812423
12912223
13212023
13010413
f2a42e23
00058913
00060493
f2d42c23
00092883
00492803
00892503
00c92583
01092603
01492683
01892703
01c92783
f1142823
f1042a23
f0a42c23
f0b42e23
f2c42023
f2d42223
f2e42423
f2f42623
f1040793
00078513
dadff0ef
fea42223
0004a883
0044a803
0084a503
00c4a583
0104a603
0144a683
0184a703
01c4a783
f1142823
f1042a23
f0a42c23
f0b42e23
f2c42023
f2d42223
f2e42423
f2f42623
f1040793
00078513
d5dff0ef
fea42023
fe442783
0a078463
fa040793
00078513
f58ff0ef
fa042883
fa442803
fa842503
fac42583
fb042603
fb442683
fb842703
fbc42783
f1142823
f1042a23
f0a42c23
f0b42e23
f2c42023
f2d42223
f2e42423
f2f42623
00092883
00492803
00892503
00c92583
01092603
01492683
01892703
01c92783
ef142823
ef042a23
eea42c23
eeb42e23
f0c42023
f0d42223
f0e42423
f0f42623
ef040713
f1040793
00070613
00078593
00090513
8d5ff0ef
fe042783
0a078463
fc040793
00078513
eacff0ef
fc042883
fc442803
fc842503
fcc42583
fd042603
fd442683
fd842703
fdc42783
ef142823
ef042a23
eea42c23
eeb42e23
f0c42023
f0d42223
f0e42423
f0f42623
0004a883
0044a803
0084a503
00c4a583
0104a603
0144a683
0184a703
01c4a783
f1142823
f1042a23
f0a42c23
f0b42e23
f2c42023
f2d42223
f2e42423
f2f42623
f1040713
ef040793
00070613
00078593
00048513
829ff0ef
f8040793
00078513
e08ff0ef
f6040793
00078513
dfcff0ef
00100793
f6f42023
fe042623
1c80006f
ef040313
f6042883
f6442803
f6842503
f6c42583
f7042603
f7442683
f7842703
f7c42783
f1142823
f1042a23
f0a42c23
f0b42e23
f2c42023
f2d42223
f2e42423
f2f42623
f6042883
f6442803
f6842503
f6c42583
f7042603
f7442683
f7842703
f7c42783
ed142823
ed042a23
eca42c23
ecb42e23
eec42023
eed42223
eee42423
eef42623
ed040713
f1040793
00070613
00078593
00030513
de8ff0ef
ef042883
ef442803
ef842503
efc42583
f0042603
f0442683
f0842703
f0c42783
f7142023
f7042223
f6a42423
f6b42623
f6c42823
f6d42a23
f6e42c23
f6f42e23
ed040313
0004a883
0044a803
0084a503
00c4a583
0104a603
0144a683
0184a703
01c4a783
ef142823
ef042a23
eea42c23
eeb42e23
f0c42023
f0d42223
f0e42423
f0f42623
0004a883
0044a803
0084a503
00c4a583
0104a603
0144a683
0184a703
01c4a783
f1142823
f1042a23
f0a42c23
f0b42e23
f2c42023
f2d42223
f2e42423
f2f42623
f1040713
ef040793
00070613
00078593
00030513
d0cff0ef
ed042883
ed442803
ed842503
edc42583
ee042603
ee442683
ee842703
eec42783
0114a023
0104a223
00a4a423
00b4a623
00c4a823
00d4aa23
00e4ac23
00f4ae23
fec42783
00178793
fef42623
fec42703
03e00793
e2e7dae3
03f00793
fef42423
3440006f
f4040313
00092883
00492803
00892503
00c92583
01092603
01492683
01892703
01c92783
ed142823
ed042a23
eca42c23
ecb42e23
eec42023
eed42223
eee42423
eef42623
0004a883
0044a803
0084a503
00c4a583
0104a603
0144a683
0184a703
01c4a783
ef142823
ef042a23
eea42c23
eeb42e23
f0c42023
f0d42223
f0e42423
f0f42623
ef040713
ed040793
00070613
00078593
00030513
d88ff0ef
f4042883
f4442803
f4842503
f4c42583
f5042603
f5442683
f5842703
f5c42783
ed142823
ed042a23
eca42c23
ecb42e23
eec42023
eed42223
eee42423
eef42623
ed040793
00078513
915ff0ef
00050793
12079063
ed040313
f8042883
f8442803
f8842503
f8c42583
f9042603
f9442683
f9842703
f9c42783
ef142823
ef042a23
eea42c23
eeb42e23
f0c42023
f0d42223
f0e42423
f0f42623
f6042883
f6442803
f6842503
f6c42583
f7042603
f7442683
f7842703
f7c42783
f1142823
f1042a23
f0a42c23
f0b42e23
f2c42023
f2d42223
f2e42423
f2f42623
f1040713
ef040793
00070613
00078593
00030513
b1cff0ef
ed042883
ed442803
ed842503
edc42583
ee042603
ee442683
ee842703
eec42783
f9142023
f9042223
f8a42423
f8b42623
f8c42823
f8d42a23
f8e42c23
f8f42e23
f4042883
f4442803
f4842503
f4c42583
f5042603
f5442683
f5842703
f5c42783
01192023
01092223
00a92423
00b92623
00c92823
00d92a23
00e92c23
00f92e23
ed040313
f6042883
f6442803
f6842503
f6c42583
f7042603
f7442683
f7842703
f7c42783
ef142823
ef042a23
eea42c23
eeb42e23
f0c42023
f0d42223
f0e42423
f0f42623
ef040793
00078593
00030513
fd4ff0ef
ed042883
ed442803
ed842503
edc42583
ee042603
ee442683
ee842703
eec42783
f7142023
f7042223
f6a42423
f6b42623
f6c42823
f6d42a23
f6e42c23
f6f42e23
ed040313
0004a883
0044a803
0084a503
00c4a583
0104a603
0144a683
0184a703
01c4a783
ef142823
ef042a23
eea42c23
eeb42e23
f0c42023
f0d42223
f0e42423
f0f42623
ef040793
00078593
00030513
f40ff0ef
ed042883
ed442803
ed842503
edc42583
ee042603
ee442683
ee842703
eec42783
0114a023
0104a223
00a4a423
00b4a623
00c4a823
00d4aa23
00e4ac23
00f4ae23
fe842783
fff78793
fef42423
fe842783
ca07dee3
f3842783
00092303
00492883
00892803
00c92503
01092583
01492603
01892683
01c92703
0067a023
0117a223
0107a423
00a7a623
00b7a823
00c7aa23
00d7ac23
00e7ae23
f3c42783
f8042303
f8442883
f8842803
f8c42503
f9042583
f9442603
f9842683
f9c42703
0067a023
0117a223
0107a423
00a7a623
00b7a823
00c7aa23
00d7ac23
00e7ae23
f3c42503
12c12083
12812403
12412483
12012903
13010113
00008067
fe010113
00812e23
00912c23
01212a23
02010413
00050493
00058913
fe042623
03c0006f
fec42783
00279793
00f487b3
0007a703
fec42783
00279793
00f907b3
0007a783
00f70663
00000793
0200006f
fec42783
00178793
fef42623
fec42703
00700793
fce7d0e3
00100793
00078513
01c12403
01812483
01412903
02010113
00008067
ea010113
14112e23
14812c23
14912a23
16010413
f0a42623
00058493
f9040793
00078513
f79fe0ef
00002797
63878793
0007a883
0047a803
0087a503
00c7a583
0107a603
0147a683
0187a703
01c7a783
f7142823
f7042a23
f6a42c23
f6b42e23
f8c42023
f8d42223
f8e42423
f8f42623
f5040793
00078513
f25fe0ef
00100793
f4f42823
4840006f
fb040313
f9042883
f9442803
f9842503
f9c42583
fa042603
fa442683
fa842703
fac42783
ef142023
ef042223
eea42423
eeb42623
eec42823
eed42a23
eee42c23
eef42e23
f7042883
f7442803
f7842503
f7c42583
f8042603
f8442683
f8842703
f8c42783
ed142023
ed042223
eca42423
ecb42623
ecc42823
ecd42a23
ece42c23
ecf42e23
ec040713
ee040793
00070613
00078593
00030513
f15fe0ef
f1040313
fb042883
fb442803
fb842503
fbc42583
fc042603
fc442683
fc842703
fcc42783
ed142023
ed042223
eca42423
ecb42623
ecc42823
ecd42a23
ece42c23
ecf42e23
ec040793
00078593
00030513
c4cff0ef
f3040313
f1042883
f1442803
f1842503
f1c42583
f2042603
f2442683
f2842703
f2c42783
ed142023
ed042223
eca42423
ecb42623
ecc42823
ecd42a23
ece42c23
ecf42e23
f1042883
f1442803
f1842503
f1c42583
f2042603
f2442683
f2842703
f2c42783
ef142023
ef042223
eea42423
eeb42623
eec42823
eed42a23
eee42c23
eef42e23
ee040713
ec040793
00070613
00078593
00030513
91cff0ef
fd040313
f3042883
f3442803
f3842503
f3c42583
f4042603
f4442683
f4842703
f4c42783
ed142023
ed042223
eca42423
ecb42623
ecc42823
ecd42a23
ece42c23
ecf42e23
0004a883
0044a803
0084a503
00c4a583
0104a603
0144a683
0184a703
01c4a783
ef142023
ef042223
eea42423
eeb42623
eec42823
eed42a23
eee42c23
eef42e23
ee040713
ec040793
00070613
00078593
00030513
f05fe0ef
fd042883
fd442803
fd842503
fdc42583
fe042603
fe442683
fe842703
fec42783
ed142023
ed042223
eca42423
ecb42623
ecc42823
ecd42a23
ece42c23
ecf42e23
ec040793
00078513
a90ff0ef
00050793
0e078263
ec040313
f1042883
f1442803
f1842503
f1c42583
f2042603
f2442683
f2842703
f2c42783
ef142023
ef042223
eea42423
eeb42623
eec42823
eed42a23
eee42c23
eef42e23
f5042883
f5442803
f5842503
f5c42583
f6042603
f6442683
f6842703
f6c42783
eb142023
eb042223
eaa42423
eab42623
eac42823
ead42a23
eae42c23
eaf42e23
ea040713
ee040793
00070613
00078593
00030513
c99fe0ef
ec042883
ec442803
ec842503
ecc42583
ed042603
ed442683
ed842703
edc42783
f9142823
f9042a23
f8a42c23
f8b42e23
fac42023
fad42223
fae42423
faf42623
1280006f
0004a883
0044a803
0084a503
00c4a583
0104a603
0144a683
0184a703
01c4a783
eb142023
eb042223
eaa42423
eab42623
eac42823
ead42a23
eae42c23
eaf42e23
f3042883
f3442803
f3842503
f3c42583
f4042603
f4442683
f4842703
f4c42783
ed142023
ed042223
eca42423
ecb42623
ecc42823
ecd42a23
ece42c23
ecf42e23
ec040713
ea040793
00070593
00078513
b09ff0ef
00050793
04078663
f0c42783
f1042303
f1442883
f1842803
f1c42503
f2042583
f2442603
f2842683
f2c42703
0067a023
0117a223
0107a423
00a7a623
00b7a823
00c7aa23
00d7ac23
00e7ae23
1240006f
f1042883
f1442803
f1842503
f1c42583
f2042603
f2442683
f2842703
f2c42783
f7142823
f7042a23
f6a42c23
f6b42e23
f8c42023
f8d42223
f8e42423
f8f42623
f9042883
f9442803
f9842503
f9c42583
fa042603
fa442683
fa842703
fac42783
eb142023
eb042223
eaa42423
eab42623
eac42823
ead42a23
eae42c23
eaf42e23
f7042883
f7442803
f7842503
f7c42583
f8042603
f8442683
f8842703
f8c42783
ed142023
ed042223
eca42423
ecb42623
ecc42823
ecd42a23
ece42c23
ecf42e23
ec040713
ea040793
00070593
00078513
9e5ff0ef
00050793
ae0784e3
f0c42783
f9042303
f9442883
f9842803
f9c42503
fa042583
fa442603
fa842683
fac42703
0067a023
0117a223
0107a423
00a7a623
00b7a823
00c7aa23
00d7ac23
00e7ae23
f0c42503
15c12083
15812403
15412483
16010113
00008067
f7010113
08112623
08812423
08912223
09010413
00050493
fab42e23
fe042623
0cc0006f
0004a883
0044a803
0084a503
00c4a583
0104a603
0144a683
0184a703
01c4a783
f9142823
f9042a23
f8a42c23
f8b42e23
fac42023
fad42223
fae42423
faf42623
00002797
f9c78793
0007a883
0047a803
0087a503
00c7a583
0107a603
0147a683
0187a703
01c7a783
f7142823
f7042a23
f6a42c23
f6b42e23
f8c42023
f8d42223
f8e42423
f8f42623
fcc40693
f7040713
f9040793
00070613
00078593
00048513
8a8ff0ef
fcc42683
fec42783
fbc42703
00f707b3
0ff6f713
00e78023
fec42783
00178793
fef42623
fec42703
00b00793
f2e7d8e3
00000013
00000013
08c12083
08812403
08412483
09010113
00008067
fe010113
00112e23
00812c23
02010413
fea42623
fec42503
821fe0ef
00050793
00078593
fec42503
ea0fe0ef
00000013
01c12083
01812403
02010113
00008067
f7010113
08112623
08812423
08912223
09010413
00050493
0004a883
0044a803
0084a503
00c4a583
0104a603
0144a683
0184a703
01c4a783
f9142823
f9042a23
f8a42c23
f8b42e23
fac42023
fad42223
fae42423
faf42623
f9040793
00078513
dd5fe0ef
00050793
0a078c63
00002517
d6c50513
f4dff0ef
fc840793
00078513
fc8fe0ef
fc842883
fcc42803
fd042503
fd442583
fd842603
fdc42683
fe042703
fe442783
f9142823
f9042a23
f8a42c23
f8b42e23
fac42023
fad42223
fae42423
faf42623
0004a883
0044a803
0084a503
00c4a583
0104a603
0144a683
0184a703
01c4a783
f7142823
f7042a23
f6a42c23
f6b42e23
f8c42023
f8d42223
f8e42423
f8f42623
f7040713
f9040793
00070613
00078593
00048513
945fe0ef
0100006f
00002517
cbc50513
e99ff0ef
0004a883
0044a803
0084a503
00c4a583
0104a603
0144a683
0184a703
01c4a783
f7142823
f7042a23
f6a42c23
f6b42e23
f8c42023
f8d42223
f8e42423
f8f42623
fbc40713
f7040793
00070593
00078513
d31ff0ef
00100793
fef42623
00b00793
fef42423
0a40006f
fe842703
00600793
00f71463
fe042623
fe842783
ff078793
008787b3
fcc7c783
02079663
fec42783
00078a63
00002517
c1c50513
df9ff0ef
0440006f
00002517
c1050513
de9ff0ef
0340006f
fe042623
fe842783
ff078793
008787b3
fcc7c783
03078793
0ff7f793
faf40da3
fbb40793
00100593
00078513
c7cfe0ef
fe842703
00600793
00f71863
00002517
bc850513
d9dff0ef
fe842783
fff78793
fef42423
fe842783
f407dee3
00000013
00000013
08c12083
08812403
08412483
09010113
00008067
f8010113
06112e23
06812c23
06912a23
08010413
00002497
c4048493
fc040793
00078513
dccfe0ef
fc042883
fc442803
fc842503
fcc42583
fd042603
fd442683
fd842703
fdc42783
0114a023
0104a223
00a4a423
00b4a623
00c4a823
00d4aa23
00e4ac23
00f4ae23
00002797
bec78793
00a00713
00e7a023
00002497
c1c48493
fc040793
00078513
d68fe0ef
fc042883
fc442803
fc842503
fcc42583
fd042603
fd442683
fd842703
fdc42783
0114a023
0104a223
00a4a423
00b4a623
00c4a823
00d4aa23
00e4ac23
00f4ae23
00002797
bc878793
00100713
00e7a023
fe042623
1600006f
fec42703
00300793
04f71a63
00002797
b8478793
00002717
b9c70713
00072303
00472883
00872803
00c72503
01072583
01472603
01872683
01c72703
0067a023
0117a223
0107a423
00a7a623
00b7a823
00c7aa23
00d7ac23
00e7ae23
00002497
b5448493
fc040313
00002797
b4878793
0007a883
0047a803
0087a503
00c7a583
0107a603
0147a683
0187a703
01c7a783
fb142023
fb042223
faa42423
fab42623
fac42823
fad42a23
fae42c23
faf42e23
00002797
ac078793
0007a883
0047a803
0087a503
00c7a583
0107a603
0147a683
0187a703
01c7a783
f9142023
f9042223
f8a42423
f8b42623
f8c42823
f8d42a23
f8e42c23
f8f42e23
f8040713
fa040793
00070613
00078593
00030513
f90fe0ef
fc042883
fc442803
fc842503
fcc42583
fd042603
fd442683
fd842703
fdc42783
0114a023
0104a223
00a4a423
00b4a623
00c4a823
00d4aa23
00e4ac23
00f4ae23
fec42783
00178793
fef42623
fec42703
00500793
e8e7dee3
00002497
a6848493
f8040313
00002797
a3c78793
0007a883
0047a803
0087a503
00c7a583
0107a603
0147a683
0187a703
01c7a783
fb142023
fb042223
faa42423
fab42623
fac42823
fad42a23
fae42c23
faf42e23
00002797
9f478793
0007a883
0047a803
0087a503
00c7a583
0107a603
0147a683
0187a703
01c7a783
fd142023
fd042223
fca42423
fcb42623
fcc42823
fcd42a23
fce42c23
fcf42e23
fc040713
fa040793
00070613
00078593
00030513
e84fe0ef
f8042883
f8442803
f8842503
f8c42583
f9042603
f9442683
f9842703
f9c42783
0114a023
0104a223
00a4a423
00b4a623
00c4a823
00d4aa23
00e4ac23
00f4ae23
00002797
99478793
0007a023
00002497
98848493
f8040793
00078513
a94fe0ef
f8042883
f8442803
f8842503
f8c42583
f9042603
f9442683
f9842703
f9c42783
0714a223
0704a423
06a4a623
06b4a823
06c4aa23
06d4ac23
06e4ae23
08f4a023
00002797
93478793
00002717
92c70713
06472303
06872883
06c72803
07072503
07472583
07872603
07c72683
08072703
0467a223
0517a423
0507a623
04a7a823
04b7aa23
04c7ac23
04d7ae23
06e7a023
00002797
8e478793
00002717
8dc70713
04472303
04872883
04c72803
05072503
05472583
05872603
05c72683
06072703
0267a223
0317a423
0307a623
02a7a823
02b7aa23
02c7ac23
02d7ae23
04e7a023
00002797
89478793
00002717
88c70713
02472303
02872883
02c72803
03072503
03472583
03872603
03c72683
04072703
0067a223
0117a423
0107a623
00a7a823
00b7aa23
00c7ac23
00d7ae23
02e7a023
00002797
84478793
0807a223
00002797
83878793
0807a423
00002797
82c78793
02000713
08e78623
00000013
07c12083
07812403
07412483
08010113
00008067
e5010113
1a112623
1a812423
1a912223
1b010413
00050793
eaf40fa3
fe042423
ee440793
00078513
8f8fe0ef
ebf44703
02f00793
78e7fa63
ebf44703
03900793
78e7e463
00001797
7c078793
ebf44703
08e78623
00001797
7b078793
0887a783
14078a63
00001797
7a078793
0807a423
00001797
79478793
00001717
78c70713
04472303
04872883
04c72803
05072503
05472583
05872603
05c72683
06072703
0667a223
0717a423
0707a623
06a7a823
06b7aa23
06c7ac23
06d7ae23
08e7a023
00001797
74478793
00001717
73c70713
02472303
02872883
02c72803
03072503
03472583
03872603
03c72683
04072703
0467a223
0517a423
0507a623
04a7a823
04b7aa23
04c7ac23
04d7ae23
06e7a023
00001797
6f478793
00001717
6ec70713
00472303
00872883
00c72803
01072503
01472583
01872603
01c72683
02072703
0267a223
0317a423
0307a623
02a7a823
02b7aa23
02c7ac23
02d7ae23
04e7a023
00001497
6a448493
e9040793
00078513
fb1fd0ef
e9042883
e9442803
e9842503
e9c42583
ea042603
ea442683
ea842703
eac42783
0114a223
0104a423
00a4a623
00b4a823
00c4aa23
00d4ac23
00e4ae23
02f4a023
ebf44783
fd078793
fef42223
00001797
64478793
0007a783
28079a63
00001497
63448493
e9040313
00001797
62878793
0047a883
0087a803
00c7a503
0107a583
0147a603
0187a683
01c7a703
0207a783
e7142823
e7042a23
e6a42c23
e6b42e23
e8c42023
e8d42223
e8e42423
e8f42623
00001797
56078793
0007a883
0047a803
0087a503
00c7a583
0107a603
0147a683
0187a703
01c7a783
e5142823
e5042a23
e4a42c23
e4b42e23
e6c42023
e6d42223
e6e42423
e6f42623
e5040713
e7040793
00070613
00078593
00030513
a30fe0ef
e9042883
e9442803
e9842503
e9c42583
ea042603
ea442683
ea842703
eac42783
0114a223
0104a423
00a4a623
00b4a823
00c4aa23
00d4ac23
00e4ae23
02f4a023
fe442783
eef42223
f0440313
ee442883
ee842803
eec42503
ef042583
ef442603
ef842683
efc42703
f0042783
e5142823
e5042a23
e4a42c23
e4b42e23
e6c42023
e6d42223
e6e42423
e6f42623
00001797
4b478793
0007a883
0047a803
0087a503
00c7a583
0107a603
0147a683
0187a703
01c7a783
e7142823
e7042a23
e6a42c23
e6b42e23
e8c42023
e8d42223
e8e42423
e8f42623
e7040713
e5040793
00070613
00078593
00030513
944fe0ef
00001497
49448493
e5040313
00001797
48878793
0047a883
0087a803
00c7a503
0107a583
0147a603
0187a683
01c7a703
0207a783
e7142823
e7042a23
e6a42c23
e6b42e23
e8c42023
e8d42223
e8e42423
e8f42623
f0442883
f0842803
f0c42503
f1042583
f1442603
f1842683
f1c42703
f2042783
e9142823
e9042a23
e8a42c23
e8b42e23
eac42023
ead42223
eae42423
eaf42623
e9040713
e7040793
00070613
00078593
00030513
da1fd0ef
e5042883
e5442803
e5842503
e5c42583
e6042603
e6442683
e6842703
e6c42783
0114a223
0104a423
00a4a623
00b4a823
00c4aa23
00d4ac23
00e4ae23
02f4a023
5300006f
00001797
3a478793
0007a703
00700793
50f70e63
00001797
35078793
0007a883
0047a803
0087a503
00c7a583
0107a603
0147a683
0187a703
01c7a783
ef142223
ef042423
eea42623
eeb42823
eec42a23
eed42c23
eee42e23
f0f42023
fe042623
0f80006f
e5040313
ee442883
ee842803
eec42503
ef042583
ef442603
ef842683
efc42703
f0042783
e7142823
e7042a23
e6a42c23
e6b42e23
e8c42023
e8d42223
e8e42423
e8f42623
00001797
27c78793
0007a883
0047a803
0087a503
00c7a583
0107a603
0147a683
0187a703
01c7a783
e9142823
e9042a23
e8a42c23
e8b42e23
eac42023
ead42223
eae42423
eaf42623
ec440693
e9040713
e7040793
00070613
00078593
00030513
b88fe0ef
e5042883
e5442803
e5842503
e5c42583
e6042603
e6442683
e6842703
e6c42783
ef142223
ef042423
eea42623
eeb42823
eec42a23
eed42c23
eee42e23
f0f42023
fec42783
00178793
fef42623
00001797
24c78793
0007a783
fec42703
eef74ee3
e5040793
00078513
b4dfd0ef
e5042883
e5442803
e5842503
e5c42583
e6042603
e6442683
e6842703
e6c42783
ed142223
ed042423
eca42623
ecb42823
ecc42a23
ecd42c23
ece42e23
eef42023
fe442783
ecf42223
f2440313
ee442883
ee842803
eec42503
ef042583
ef442603
ef842683
efc42703
f0042783
e5142823
e5042a23
e4a42c23
e4b42e23
e6c42023
e6d42223
e6e42423
e6f42623
ec442883
ec842803
ecc42503
ed042583
ed442603
ed842683
edc42703
ee042783
e7142823
e7042a23
e6a42c23
e6b42e23
e8c42023
e8d42223
e8e42423
e8f42623
e7040713
e5040793
00070613
00078593
00030513
df9fd0ef
00001497
14848493
e5040313
00001797
13c78793
0047a883
0087a803
00c7a503
0107a583
0147a603
0187a683
01c7a703
0207a783
e7142823
e7042a23
e6a42c23
e6b42e23
e8c42023
e8d42223
e8e42423
e8f42623
f2442883
f2842803
f2c42503
f3042583
f3442603
f3842683
f3c42703
f4042783
e9142823
e9042a23
e8a42c23
e8b42e23
eac42023
ead42223
eae42423
eaf42623
e9040713
e7040793
00070613
00078593
00030513
a55fd0ef
e5042883
e5442803
e5842503
e5c42583
e6042603
e6442683
e6842703
e6c42783
0114a223
0104a423
00a4a623
00b4a823
00c4aa23
00d4ac23
00e4ae23
02f4a023
00001797
05c78793
0007a783
00178713
00001797
04c78793
00e7a023
1c80006f
ebf44703
02e00793
02f71c63
00001797
03078793
0007a783
1a079863
00001797
02078793
00100713
00e7a023
00001797
01078793
02e00713
08e78623
18c0006f
ebf44703
00d00793
16f71463
00001797
ff078793
03b00713
08e78623
00001797
fe078793
00001717
fd870713
04472303
04872883
04c72803
05072503
05472583
05872603
05c72683
06072703
0667a223
0717a423
0707a623
06a7a823
06b7aa23
06c7ac23
06d7ae23
08e7a023
00001797
f9078793
00001717
f8870713
02472303
02872883
02c72803
03072503
03472583
03872603
03c72683
04072703
0467a223
0517a423
0507a623
04a7a823
04b7aa23
04c7ac23
04d7ae23
06e7a023
00001797
f4078793
00001717
f3870713
00472303
00872883
00c72803
01072503
01472583
01872603
01c72683
02072703
0267a223
0317a423
0307a623
02a7a823
02b7aa23
02c7ac23
02d7ae23
04e7a023
00001497
ef048493
e5040793
00078513
ffcfd0ef
e5042883
e5442803
e5842503
e5c42583
e6042603
e6442683
e6842703
e6c42783
0114a223
0104a423
00a4a623
00b4a823
00c4aa23
00d4ac23
00e4ae23
02f4a023
00001797
e9c78793
0007a023
01c0006f
ebf44703
07200793
00f71863
9acff0ef
0080006f
00000013
ebf44703
02b00793
02f70463
ebf44703
02d00793
00f70e63
ebf44703
02a00793
00f70863
ebf44703
02f00793
60f71a63
00001797
e4478793
ebf44703
08e78623
ebf44703
02b00793
0ef71c63
00001497
e2848493
e5040313
00001797
e1c78793
0047a883
0087a803
00c7a503
0107a583
0147a603
0187a683
01c7a703
0207a783
e7142823
e7042a23
e6a42c23
e6b42e23
e8c42023
e8d42223
e8e42423
e8f42623
00001797
dd478793
0247a883
0287a803
02c7a503
0307a583
0347a603
0387a683
03c7a703
0407a783
e9142823
e9042a23
e8a42c23
e8b42e23
eac42023
ead42223
eae42423
eaf42623
e9040713
e7040793
00070613
00078593
00030513
f2cfd0ef
e5042883
e5442803
e5842503
e5c42583
e6042603
e6442683
e6842703
e6c42783
0114a223
0104a423
00a4a623
00b4a823
00c4aa23
00d4ac23
00e4ae23
02f4a023
ebf44703
02d00793
0ef71c63
00001497
d2848493
e5040313
00001797
d1c78793
0247a883
0287a803
02c7a503
0307a583
0347a603
0387a683
03c7a703
0407a783
e7142823
e7042a23
e6a42c23
e6b42e23
e8c42023
e8d42223
e8e42423
e8f42623
00001797
cd478793
0047a883
0087a803
00c7a503
0107a583
0147a603
0187a683
01c7a703
0207a783
e9142823
e9042a23
e8a42c23
e8b42e23
eac42023
ead42223
eae42423
eaf42623
e9040713
e7040793
00070613
00078593
00030513
fa8fd0ef
e5042883
e5442803
e5842503
e5c42583
e6042603
e6442683
e6842703
e6c42783
0114a223
0104a423
00a4a623
00b4a823
00c4aa23
00d4ac23
00e4ae23
02f4a023
ebf44703
02a00793
1af71063
f4440313
00001797
c2478793
0047a883
0087a803
00c7a503
0107a583
0147a603
0187a683
01c7a703
0207a783
e5142823
e5042a23
e4a42c23
e4b42e23
e6c42023
e6d42223
e6e42423
e6f42623
00001797
bdc78793
0247a883
0287a803
02c7a503
0307a583
0347a603
0387a683
03c7a703
0407a783
e7142823
e7042a23
e6a42c23
e6b42e23
e8c42023
e8d42223
e8e42423
e8f42623
e7040713
e5040793
00070613
00078593
00030513
82dfd0ef
00001497
b7c48493
e5040313
f4442883
f4842803
f4c42503
f5042583
f5442603
f5842683
f5c42703
f6042783
e7142823
e7042a23
e6a42c23
e6b42e23
e8c42023
e8d42223
e8e42423
e8f42623
00001797
af078793
0007a883
0047a803
0087a503
00c7a583
0107a603
0147a683
0187a703
01c7a783
e9142823
e9042a23
e8a42c23
e8b42e23
eac42023
ead42223
eae42423
eaf42623
ee440693
e9040713
e7040793
00070613
00078593
00030513
bbdfd0ef
e5042883
e5442803
e5842503
e5c42583
e6042603
e6442683
e6842703
e6c42783
0114a223
0104a423
00a4a623
00b4a823
00c4aa23
00d4ac23
00e4ae23
02f4a023
ebf44703
02f00793
1af71063
f6440313
00001797
a7c78793
0247a883
0287a803
02c7a503
0307a583
0347a603
0387a683
03c7a703
0407a783
e5142823
e5042a23
e4a42c23
e4b42e23
e6c42023
e6d42223
e6e42423
e6f42623
00001797
a3478793
0047a883
0087a803
00c7a503
0107a583
0147a603
0187a683
01c7a703
0207a783
e7142823
e7042a23
e6a42c23
e6b42e23
e8c42023
e8d42223
e8e42423
e8f42623
ee440693
e7040713
e5040793
00070613
00078593
00030513
ac1fd0ef
00001497
9d048493
e5040313
f6442883
f6842803
f6c42503
f7042583
f7442603
f7842683
f7c42703
f8042783
e7142823
e7042a23
e6a42c23
e6b42e23
e8c42023
e8d42223
e8e42423
e8f42623
00001797
94478793
0007a883
0047a803
0087a503
00c7a583
0107a603
0147a683
0187a703
01c7a783
e9142823
e9042a23
e8a42c23
e8b42e23
eac42023
ead42223
eae42423
eaf42623
e9040713
e7040793
00070613
00078593
00030513
dd4fd0ef
e5042883
e5442803
e5842503
e5c42583
e6042603
e6442683
e6842703
e6c42783
0114a223
0104a423
00a4a623
00b4a823
00c4aa23
00d4ac23
00e4ae23
02f4a023
00001797
8e478793
00001717
8dc70713
04472303
04872883
04c72803
05072503
05472583
05872603
05c72683
06072703
0267a223
0317a423
0307a623
02a7a823
02b7aa23
02c7ac23
02d7ae23
04e7a023
00001797
89478793
00001717
88c70713
06472303
06872883
06c72803
07072503
07472583
07872603
07c72683
08072703
0467a223
0517a423
0507a623
04a7a823
04b7aa23
04c7ac23
04d7ae23
06e7a023
00001797
84478793
00100713
08e7a423
ebf44703
07300793
14f71e63
f8440313
00001797
82478793
0047a883
0087a803
00c7a503
0107a583
0147a603
0187a683
01c7a703
0207a783
e5142823
e5042a23
e4a42c23
e4b42e23
e6c42023
e6d42223
e6e42423
e6f42623
00000797
79c78793
0007a883
0047a803
0087a503
00c7a583
0107a603
0147a683
0187a703
01c7a783
e7142823
e7042a23
e6a42c23
e6b42e23
e8c42023
e8d42223
e8e42423
e8f42623
e7040713
e5040793
00070613
00078593
00030513
c2cfd0ef
00000497
77c48493
e5040313
f8442883
f8842803
f8c42503
f9042583
f9442603
f9842683
f9c42703
fa042783
e7142823
e7042a23
e6a42c23
e6b42e23
e8c42023
e8d42223
e8e42423
e8f42623
e7040793
00078593
00030513
8a4fe0ef
e5042883
e5442803
e5842503
e5c42583
e6042603
e6442683
e6842703
e6c42783
0114a223
0104a423
00a4a623
00b4a823
00c4aa23
00d4ac23
00e4ae23
02f4a023
00000797
6e078793
00100713
08e7a423
00000797
6d078793
0847a783
02078463
ebf44703
00d00793
00f70e63
ebf44703
00a00793
00f70863
00000797
6a878793
0807a223
00000797
69c78793
0047a883
0087a803
00c7a503
0107a583
0147a603
0187a683
01c7a703
0207a783
ef142223
ef042423
eea42623
eeb42823
eec42a23
eed42c23
eee42e23
f0f42023
ee442883
ee842803
eec42503
ef042583
ef442603
ef842683
efc42703
f0042783
e5142823
e5042a23
e4a42c23
e4b42e23
e6c42023
e6d42223
e6e42423
e6f42623
e5040793
00078513
d14fd0ef
00050793
0e078663
fa440793
00078513
f15fc0ef
e5040313
fa442883
fa842803
fac42503
fb042583
fb442603
fb842683
fbc42703
fc042783
e7142823
e7042a23
e6a42c23
e6b42e23
e8c42023
e8d42223
e8e42423
e8f42623
ee442883
ee842803
eec42503
ef042583
ef442603
ef842683
efc42703
f0042783
e9142823
e9042a23
e8a42c23
e8b42e23
eac42023
ead42223
eae42423
eaf42623
e9040713
e7040793
00070613
00078593
00030513
88cfd0ef
e5042883
e5442803
e5842503
e5c42583
e6042603
e6442683
e6842703
e6c42783
ef142223
ef042423
eea42623
eeb42823
eec42a23
eed42c23
eee42e23
f0f42023
fc440313
ee442883
ee842803
eec42503
ef042583
ef442603
ef842683
efc42703
f0042783
e5142823
e5042a23
e4a42c23
e4b42e23
e6c42023
e6d42223
e6e42423
e6f42623
00000797
4b478793
0007a883
0047a803
0087a503
00c7a583
0107a603
0147a683
0187a703
01c7a783
e7142823
e7042a23
e6a42c23
e6b42e23
e8c42023
e8d42223
e8e42423
e8f42623
e7040713
e5040793
00070613
00078593
00030513
fa9fc0ef
fc442883
fc842803
fcc42503
fd042583
fd442603
fd842683
fdc42703
fe042783
e5142823
e5042a23
e4a42c23
e4b42e23
e6c42023
e6d42223
e6e42423
e6f42623
e5040793
00078513
b34fd0ef
00050793
06079463
00000797
42078793
00100713
08e7a223
00000497
41048493
e5040793
00078513
d1dfc0ef
e5042883
e5442803
e5842503
e5c42583
e6042603
e6442683
e6842703
e6c42783
0114a223
0104a423
00a4a623
00b4a823
00c4aa23
00d4ac23
00e4ae23
02f4a023
00000013
1ac12083
1a812403
1a412483
1b010113
00008067
fd010113
02112623
02812423
03010413
00000797
31078793
0007a023
eb4fe0ef
00000517
24050513
c10fe0ef
00000517
24850513
c04fe0ef
00000517
24850513
bf8fe0ef
00000517
27c50513
becfe0ef
00000797
35478793
0647a883
0687a803
06c7a503
0707a583
0747a603
0787a683
07c7a703
0807a783
fd142823
fd042a23
fca42c23
fcb42e23
fec42023
fed42223
fee42423
fef42623
fd040793
00078513
bd8fe0ef
00000517
22450513
b8cfe0ef
00000517
21c50513
b80fe0ef
00000797
2e878793
0447a883
0487a803
04c7a503
0507a583
0547a603
0587a683
05c7a703
0607a783
fd142823
fd042a23
fca42c23
fcb42e23
fec42023
fed42223
fee42423
fef42623
fd040793
00078513
b6cfe0ef
00000517
1b850513
b20fe0ef
00000517
1b850513
b14fe0ef
00000797
27c78793
0247a883
0287a803
02c7a503
0307a583
0347a603
0387a683
03c7a703
0407a783
fd142823
fd042a23
fca42c23
fcb42e23
fec42023
fed42223
fee42423
fef42623
fd040793
00078513
b00fe0ef
00000517
14c50513
ab4fe0ef
00000517
15450513
aa8fe0ef
00000797
21078793
0047a883
0087a803
00c7a503
0107a583
0147a603
0187a683
01c7a703
0207a783
fd142823
fd042a23
fca42c23
fcb42e23
fec42023
fed42223
fee42423
fef42623
fd040793
00078513
a94fe0ef
00000517
0e050513
a48fe0ef
00000797
1b078793
0847a783
00078863
00000517
0ec50513
a2cfe0ef
00000517
0b850513
a20fe0ef
00000517
0f450513
a14fe0ef
00100593
00000517
20450513
8cdfc0ef
99dfc0ef
00050793
00078513
95dfe0ef
de5ff06f
ffff0000
0000002d
00000020
00000030
0000002e
2d524159
636c6143
74616c75
0a0d726f
00000000
325b201b
5b201b4a
0000483b
335b201b
36343b30
4159206d
72502d52
7365636f
20726f73
6c707041
74616369
206e6f69
6f6d6544
5052203a
6143204e
6c75636c
726f7461
305b201b
000d0a6d
203a5409
00000000
00000d0a
203a5a09
00000000
203a5909
00000000
5b201b09
343b3733
3a586d34
5b201b20
00006d30
335b201b
31343b37
5241576d
474e494e
764f203a
6c667265
201b776f
006d305b
7473614c
79654b20
0000203a
80000000
