00007137
00007437
00003517
54c50513
00050067
fd010113
02812623
03010413
fca42e23
fcb42c23
0a40006f
00004797
89078793
0007a783
0007c783
fef407a3
fef44783
0047d793
fef40723
fef44783
00f7f793
fef406a3
fed44783
00178793
0ff7f793
00f7f793
fef40623
fec44703
fee44783
00f71463
0540006f
00004797
84078793
0007a703
fed44783
02078793
00f707b3
fdc42703
00074703
00e78023
00004797
81c78793
0007a783
fec44703
00e78023
fdc42783
00178793
fcf42e23
fd842783
fff78793
fcf42c23
fd842783
f4079ee3
00000013
00000013
02c12403
03010113
00008067
fe010113
00812e23
02010413
00003797
7c878793
0007a783
0017c783
fef407a3
fef44783
00f7f793
fef407a3
fef44703
00003797
7a878793
0007a783
fcf708e3
00003797
79478793
0007a703
00003797
78c78793
0007a783
01078793
00f707b3
0007c783
fef40723
00003797
77078793
0007a783
00178793
00f7f713
00003797
75c78793
00e7a023
fee44783
00078513
01c12403
02010113
00008067
fd010113
02812623
03010413
fca42e23
fe042623
01c0006f
fec42783
00178793
fef42623
fdc42783
00178793
fcf42e23
fdc42783
0007c783
fe0790e3
fec42783
00078513
02c12403
03010113
00008067
fb010113
04812623
05010413
faa42e23
fe042623
0240006f
fec42783
00279793
ff078793
008787b3
fc07ae23
fec42783
00178793
fef42623
fec42703
00700793
fce7dce3
fbc42783
fcc42303
fd042883
fd442803
fd842503
fdc42583
fe042603
fe442683
fe842703
0067a023
0117a223
0107a423
00a7a623
00b7a823
00c7aa23
00d7ac23
00e7ae23
fbc42503
04c12403
05010113
00008067
fb010113
04112623
04812423
04912223
05212023
05010413
faa42e23
00058493
00060913
fcc40793
00078513
f3dff0ef
fe042623
0dc0006f
fec42783
00279793
00f487b3
0007a703
fec42783
00279793
00f907b3
0007a783
00f70733
fec42783
00279793
ff078793
008787b3
fdc7a783
00f70733
fec42783
00279793
ff078793
008787b3
fce7ae23
fec42783
00279793
ff078793
008787b3
fdc7a703
ffff07b7
00f777b3
06078063
fec42783
00279793
ff078793
008787b3
fdc7a703
ffff07b7
fff7c793
00f77733
fec42783
00279793
ff078793
008787b3
fce7ae23
fec42703
00700793
02f70063
fec42783
00178793
00279793
ff078793
008787b3
00100713
fce7ae23
fec42783
00178793
fef42623
fec42703
00700793
f2e7d0e3
fbc42783
fcc42303
fd042883
fd442803
fd842503
fdc42583
fe042603
fe442683
fe842703
0067a023
0117a223
0107a423
00a7a623
00b7a823
00c7aa23
00d7ac23
00e7ae23
fbc42503
04c12083
04812403
04412483
04012903
05010113
00008067
fb010113
04112623
04812423
04912223
05212023
05010413
faa42e23
00058493
00060913
fcc40793
00078513
dc1ff0ef
fe042623
0dc0006f
fec42783
00279793
00f487b3
0007a703
fec42783
00279793
00f907b3
0007a783
40f70733
fec42783
00279793
ff078793
008787b3
fdc7a783
40f70733
fec42783
00279793
ff078793
008787b3
fce7ae23
fec42783
00279793
ff078793
008787b3
fdc7a703
ffff07b7
00f777b3
06078063
fec42783
00279793
ff078793
008787b3
fdc7a703
ffff07b7
fff7c793
00f77733
fec42783
00279793
ff078793
008787b3
fce7ae23
fec42703
00700793
02f70063
fec42783
00178793
00279793
ff078793
008787b3
00100713
fce7ae23
fec42783
00178793
fef42623
fec42703
00700793
f2e7d0e3
fbc42783
fcc42303
fd042883
fd442803
fd842503
fdc42583
fe042603
fe442683
fe842703
0067a023
0117a223
0107a423
00a7a623
00b7a823
00c7aa23
00d7ac23
00e7ae23
fbc42503
04c12083
04812403
04412483
04012903
05010113
00008067
f5010113
0a112623
0a812423
0a912223
0b212023
0b010413
faa42e23
00058493
00060913
fcc40793
00078513
c45ff0ef
fe042623
1bc0006f
fec42783
41f7d713
00f77713
00f707b3
4047d793
00279793
00f907b3
0007a783
fec42703
00f77713
00100693
00e69733
00e7f7b3
0e078063
f9040313
fcc42883
fd042803
fd442503
fd842583
fdc42603
fe042683
fe442703
fe842783
f7142823
f7042a23
f6a42c23
f6b42e23
f8c42023
f8d42223
f8e42423
f8f42623
0004a883
0044a803
0084a503
00c4a583
0104a603
0144a683
0184a703
01c4a783
f5142823
f5042a23
f4a42c23
f4b42e23
f6c42023
f6d42223
f6e42423
f6f42623
f5040713
f7040793
00070613
00078593
00030513
c01ff0ef
f9042883
f9442803
f9842503
f9c42583
fa042603
fa442683
fa842703
fac42783
fd142623
fd042823
fca42a23
fcb42c23
fcc42e23
fed42023
fee42223
fef42423
0004a883
0044a803
0084a503
00c4a583
0104a603
0144a683
0184a703
01c4a783
f5142823
f5042a23
f4a42c23
f4b42e23
f6c42023
f6d42223
f6e42423
f6f42623
0004a883
0044a803
0084a503
00c4a583
0104a603
0144a683
0184a703
01c4a783
f7142823
f7042a23
f6a42c23
f6b42e23
f8c42023
f8d42223
f8e42423
f8f42623
f7040713
f5040793
00070613
00078593
00048513
b29ff0ef
fec42783
00178793
fef42623
fec42703
07f00793
e4e7d0e3
fbc42783
fcc42303
fd042883
fd442803
fd842503
fdc42583
fe042603
fe442683
fe842703
0067a023
0117a223
0107a423
00a7a623
00b7a823
00c7aa23
00d7ac23
00e7ae23
fbc42503
0ac12083
0a812403
0a412483
0a012903
0b010113
00008067
ff010113
00812623
00912423
01010413
00050493
01c4a783
00179713
ffff07b7
00f777b3
00078513
00c12403
00812483
01010113
00008067
fb010113
04812623
04912423
05010413
faa42e23
00058493
0004a883
0044a803
0084a503
00c4a583
0104a603
0144a683
0184a703
01c4a783
fd142623
fd042823
fca42a23
fcb42c23
fcc42e23
fed42023
fee42223
fef42423
fe042623
0ec0006f
fec42783
00279793
ff078793
008787b3
fdc7a783
0017d713
fec42783
00279793
ff078793
008787b3
fce7ae23
fec42703
00700793
04f70e63
fec42783
00279793
ff078793
008787b3
fdc7a703
fec42783
00178793
00279793
ff078793
008787b3
fdc7a783
00f79693
000107b7
fff78793
00f6f7b3
00f76733
fec42783
00279793
ff078793
008787b3
fce7ae23
0500006f
fec42783
00279793
ff078793
008787b3
fdc7a703
fec42783
00279793
ff078793
008787b3
fdc7a783
00179693
000087b7
00f6f7b3
00f76733
fec42783
00279793
ff078793
008787b3
fce7ae23
fec42783
00178793
fef42623
fec42703
00700793
f0e7d8e3
fbc42783
fcc42303
fd042883
fd442803
fd842503
fdc42583
fe042603
fe442683
fe842703
0067a023
0117a223
0107a423
00a7a623
00b7a823
00c7aa23
00d7ac23
00e7ae23
fbc42503
04c12403
04812483
05010113
00008067
ed010113
12112623
12812423
12912223
13212023
13010413
f2a42e23
00058913
00060493
f2d42c23
00092883
00492803
00892503
00c92583
01092603
01492683
01892703
01c92783
f1142823
f1042a23
f0a42c23
f0b42e23
f2c42023
f2d42223
f2e42423
f2f42623
f1040793
00078513
dadff0ef
fea42223
0004a883
0044a803
0084a503
00c4a583
0104a603
0144a683
0184a703
01c4a783
f1142823
f1042a23
f0a42c23
f0b42e23
f2c42023
f2d42223
f2e42423
f2f42623
f1040793
00078513
d5dff0ef
fea42023
fe442783
0a078463
fa040793
00078513
f58ff0ef
fa042883
fa442803
fa842503
fac42583
fb042603
fb442683
fb842703
fbc42783
f1142823
f1042a23
f0a42c23
f0b42e23
f2c42023
f2d42223
f2e42423
f2f42623
00092883
00492803
00892503
00c92583
01092603
01492683
01892703
01c92783
ef142823
ef042a23
eea42c23
eeb42e23
f0c42023
f0d42223
f0e42423
f0f42623
ef040713
f1040793
00070613
00078593
00090513
8d5ff0ef
fe042783
0a078463
fc040793
00078513
eacff0ef
fc042883
fc442803
fc842503
fcc42583
fd042603
fd442683
fd842703
fdc42783
ef142823
ef042a23
eea42c23
eeb42e23
f0c42023
f0d42223
f0e42423
f0f42623
0004a883
0044a803
0084a503
00c4a583
0104a603
0144a683
0184a703
01c4a783
f1142823
f1042a23
f0a42c23
f0b42e23
f2c42023
f2d42223
f2e42423
f2f42623
f1040713
ef040793
00070613
00078593
00048513
829ff0ef
f8040793
00078513
e08ff0ef
f6040793
00078513
dfcff0ef
00100793
f6f42023
fe042623
1c80006f
ef040313
f6042883
f6442803
f6842503
f6c42583
f7042603
f7442683
f7842703
f7c42783
f1142823
f1042a23
f0a42c23
f0b42e23
f2c42023
f2d42223
f2e42423
f2f42623
f6042883
f6442803
f6842503
f6c42583
f7042603
f7442683
f7842703
f7c42783
ed142823
ed042a23
eca42c23
ecb42e23
eec42023
eed42223
eee42423
eef42623
ed040713
f1040793
00070613
00078593
00030513
de8ff0ef
ef042883
ef442803
ef842503
efc42583
f0042603
f0442683
f0842703
f0c42783
f7142023
f7042223
f6a42423
f6b42623
f6c42823
f6d42a23
f6e42c23
f6f42e23
ed040313
0004a883
0044a803
0084a503
00c4a583
0104a603
0144a683
0184a703
01c4a783
ef142823
ef042a23
eea42c23
eeb42e23
f0c42023
f0d42223
f0e42423
f0f42623
0004a883
0044a803
0084a503
00c4a583
0104a603
0144a683
0184a703
01c4a783
f1142823
f1042a23
f0a42c23
f0b42e23
f2c42023
f2d42223
f2e42423
f2f42623
f1040713
ef040793
00070613
00078593
00030513
d0cff0ef
ed042883
ed442803
ed842503
edc42583
ee042603
ee442683
ee842703
eec42783
0114a023
0104a223
00a4a423
00b4a623
00c4a823
00d4aa23
00e4ac23
00f4ae23
fec42783
00178793
fef42623
fec42703
03e00793
e2e7dae3
03f00793
fef42423
3440006f
f4040313
00092883
00492803
00892503
00c92583
01092603
01492683
01892703
01c92783
ed142823
ed042a23
eca42c23
ecb42e23
eec42023
eed42223
eee42423
eef42623
0004a883
0044a803
0084a503
00c4a583
0104a603
0144a683
0184a703
01c4a783
ef142823
ef042a23
eea42c23
eeb42e23
f0c42023
f0d42223
f0e42423
f0f42623
ef040713
ed040793
00070613
00078593
00030513
d88ff0ef
f4042883
f4442803
f4842503
f4c42583
f5042603
f5442683
f5842703
f5c42783
ed142823
ed042a23
eca42c23
ecb42e23
eec42023
eed42223
eee42423
eef42623
ed040793
00078513
915ff0ef
00050793
12079063
ed040313
f8042883
f8442803
f8842503
f8c42583
f9042603
f9442683
f9842703
f9c42783
ef142823
ef042a23
eea42c23
eeb42e23
f0c42023
f0d42223
f0e42423
f0f42623
f6042883
f6442803
f6842503
f6c42583
f7042603
f7442683
f7842703
f7c42783
f1142823
f1042a23
f0a42c23
f0b42e23
f2c42023
f2d42223
f2e42423
f2f42623
f1040713
ef040793
00070613
00078593
00030513
b1cff0ef
ed042883
ed442803
ed842503
edc42583
ee042603
ee442683
ee842703
eec42783
f9142023
f9042223
f8a42423
f8b42623
f8c42823
f8d42a23
f8e42c23
f8f42e23
f4042883
f4442803
f4842503
f4c42583
f5042603
f5442683
f5842703
f5c42783
01192023
01092223
00a92423
00b92623
00c92823
00d92a23
00e92c23
00f92e23
ed040313
f6042883
f6442803
f6842503
f6c42583
f7042603
f7442683
f7842703
f7c42783
ef142823
ef042a23
eea42c23
eeb42e23
f0c42023
f0d42223
f0e42423
f0f42623
ef040793
00078593
00030513
fd4ff0ef
ed042883
ed442803
ed842503
edc42583
ee042603
ee442683
ee842703
eec42783
f7142023
f7042223
f6a42423
f6b42623
f6c42823
f6d42a23
f6e42c23
f6f42e23
ed040313
0004a883
0044a803
0084a503
00c4a583
0104a603
0144a683
0184a703
01c4a783
ef142823
ef042a23
eea42c23
eeb42e23
f0c42023
f0d42223
f0e42423
f0f42623
ef040793
00078593
00030513
f40ff0ef
ed042883
ed442803
ed842503
edc42583
ee042603
ee442683
ee842703
eec42783
0114a023
0104a223
00a4a423
00b4a623
00c4a823
00d4aa23
00e4ac23
00f4ae23
fe842783
fff78793
fef42423
fe842783
ca07dee3
f3842783
00092303
00492883
00892803
00c92503
01092583
01492603
01892683
01c92703
0067a023
0117a223
0107a423
00a7a623
00b7a823
00c7aa23
00d7ac23
00e7ae23
f3c42783
f8042303
f8442883
f8842803
f8c42503
f9042583
f9442603
f9842683
f9c42703
0067a023
0117a223
0107a423
00a7a623
00b7a823
00c7aa23
00d7ac23
00e7ae23
f3c42503
12c12083
12812403
12412483
12012903
13010113
00008067
fe010113
00812e23
00912c23
01212a23
02010413
00050493
00058913
fe042623
03c0006f
fec42783
00279793
00f487b3
0007a703
fec42783
00279793
00f907b3
0007a783
00f70663
00000793
0200006f
fec42783
00178793
fef42623
fec42703
00700793
fce7d0e3
00100793
00078513
01c12403
01812483
01412903
02010113
00008067
ea010113
14112e23
14812c23
14912a23
16010413
f0a42623
00058493
f9040793
00078513
f79fe0ef
00002797
6c478793
0007a883
0047a803
0087a503
00c7a583
0107a603
0147a683
0187a703
01c7a783
f7142823
f7042a23
f6a42c23
f6b42e23
f8c42023
f8d42223
f8e42423
f8f42623
f5040793
00078513
f25fe0ef
00100793
f4f42823
4840006f
fb040313
f9042883
f9442803
f9842503
f9c42583
fa042603
fa442683
fa842703
fac42783
ef142023
ef042223
eea42423
eeb42623
eec42823
eed42a23
eee42c23
eef42e23
f7042883
f7442803
f7842503
f7c42583
f8042603
f8442683
f8842703
f8c42783
ed142023
ed042223
eca42423
ecb42623
ecc42823
ecd42a23
ece42c23
ecf42e23
ec040713
ee040793
00070613
00078593
00030513
f15fe0ef
f1040313
fb042883
fb442803
fb842503
fbc42583
fc042603
fc442683
fc842703
fcc42783
ed142023
ed042223
eca42423
ecb42623
ecc42823
ecd42a23
ece42c23
ecf42e23
ec040793
00078593
00030513
c4cff0ef
f3040313
f1042883
f1442803
f1842503
f1c42583
f2042603
f2442683
f2842703
f2c42783
ed142023
ed042223
eca42423
ecb42623
ecc42823
ecd42a23
ece42c23
ecf42e23
f1042883
f1442803
f1842503
f1c42583
f2042603
f2442683
f2842703
f2c42783
ef142023
ef042223
eea42423
eeb42623
eec42823
eed42a23
eee42c23
eef42e23
ee040713
ec040793
00070613
00078593
00030513
91cff0ef
fd040313
f3042883
f3442803
f3842503
f3c42583
f4042603
f4442683
f4842703
f4c42783
ed142023
ed042223
eca42423
ecb42623
ecc42823
ecd42a23
ece42c23
ecf42e23
0004a883
0044a803
0084a503
00c4a583
0104a603
0144a683
0184a703
01c4a783
ef142023
ef042223
eea42423
eeb42623
eec42823
eed42a23
eee42c23
eef42e23
ee040713
ec040793
00070613
00078593
00030513
f05fe0ef
fd042883
fd442803
fd842503
fdc42583
fe042603
fe442683
fe842703
fec42783
ed142023
ed042223
eca42423
ecb42623
ecc42823
ecd42a23
ece42c23
ecf42e23
ec040793
00078513
a90ff0ef
00050793
0e078263
ec040313
f1042883
f1442803
f1842503
f1c42583
f2042603
f2442683
f2842703
f2c42783
ef142023
ef042223
eea42423
eeb42623
eec42823
eed42a23
eee42c23
eef42e23
f5042883
f5442803
f5842503
f5c42583
f6042603
f6442683
f6842703
f6c42783
eb142023
eb042223
eaa42423
eab42623
eac42823
ead42a23
eae42c23
eaf42e23
ea040713
ee040793
00070613
00078593
00030513
c99fe0ef
ec042883
ec442803
ec842503
ecc42583
ed042603
ed442683
ed842703
edc42783
f9142823
f9042a23
f8a42c23
f8b42e23
fac42023
fad42223
fae42423
faf42623
1280006f
0004a883
0044a803
0084a503
00c4a583
0104a603
0144a683
0184a703
01c4a783
eb142023
eb042223
eaa42423
eab42623
eac42823
ead42a23
eae42c23
eaf42e23
f3042883
f3442803
f3842503
f3c42583
f4042603
f4442683
f4842703
f4c42783
ed142023
ed042223
eca42423
ecb42623
ecc42823
ecd42a23
ece42c23
ecf42e23
ec040713
ea040793
00070593
00078513
b09ff0ef
00050793
04078663
f0c42783
f1042303
f1442883
f1842803
f1c42503
f2042583
f2442603
f2842683
f2c42703
0067a023
0117a223
0107a423
00a7a623
00b7a823
00c7aa23
00d7ac23
00e7ae23
1240006f
f1042883
f1442803
f1842503
f1c42583
f2042603
f2442683
f2842703
f2c42783
f7142823
f7042a23
f6a42c23
f6b42e23
f8c42023
f8d42223
f8e42423
f8f42623
f9042883
f9442803
f9842503
f9c42583
fa042603
fa442683
fa842703
fac42783
eb142023
eb042223
eaa42423
eab42623
eac42823
ead42a23
eae42c23
eaf42e23
f7042883
f7442803
f7842503
f7c42583
f8042603
f8442683
f8842703
f8c42783
ed142023
ed042223
eca42423
ecb42623
ecc42823
ecd42a23
ece42c23
ecf42e23
ec040713
ea040793
00070593
00078513
9e5ff0ef
00050793
ae0784e3
f0c42783
f9042303
f9442883
f9842803
f9c42503
fa042583
fa442603
fa842683
fac42703
0067a023
0117a223
0107a423
00a7a623
00b7a823
00c7aa23
00d7ac23
00e7ae23
f0c42503
15c12083
15812403
15412483
16010113
00008067
f7010113
08112623
08812423
08912223
09010413
00050493
fab42e23
fe042623
0cc0006f
0004a883
0044a803
0084a503
00c4a583
0104a603
0144a683
0184a703
01c4a783
f9142823
f9042a23
f8a42c23
f8b42e23
fac42023
fad42223
fae42423
faf42623
00002797
02878793
0007a883
0047a803
0087a503
00c7a583
0107a603
0147a683
0187a703
01c7a783
f7142823
f7042a23
f6a42c23
f6b42e23
f8c42023
f8d42223
f8e42423
f8f42623
fcc40693
f7040713
f9040793
00070613
00078593
00048513
8a8ff0ef
fcc42683
fec42783
fbc42703
00f707b3
0ff6f713
00e78023
fec42783
00178793
fef42623
fec42703
00b00793
f2e7d8e3
00000013
00000013
08c12083
08812403
08412483
09010113
00008067
fe010113
00112e23
00812c23
02010413
fea42623
fec42503
821fe0ef
00050793
00078593
fec42503
ea0fe0ef
00000013
01c12083
01812403
02010113
00008067
f6010113
08112e23
08812c23
08912a23
0a010413
00050493
fab42623
0004a883
0044a803
0084a503
00c4a583
0104a603
0144a683
0184a703
01c4a783
f9142023
f9042223
f8a42423
f8b42623
f8c42823
f8d42a23
f8e42c23
f8f42e23
f8040793
00078513
dd1fe0ef
00050793
0c078063
fac42783
00178713
fae42623
02d00713
00e78023
fc840793
00078513
fbcfe0ef
fc842883
fcc42803
fd042503
fd442583
fd842603
fdc42683
fe042703
fe442783
f9142023
f9042223
f8a42423
f8b42623
f8c42823
f8d42a23
f8e42c23
f8f42e23
0004a883
0044a803
0084a503
00c4a583
0104a603
0144a683
0184a703
01c4a783
f7142023
f7042223
f6a42423
f6b42623
f6c42823
f6d42a23
f6e42c23
f6f42e23
f6040713
f8040793
00070613
00078593
00048513
939fe0ef
0180006f
fac42783
00178713
fae42623
02000713
00e78023
0004a883
0044a803
0084a503
00c4a583
0104a603
0144a683
0184a703
01c4a783
f7142023
f7042223
f6a42423
f6b42623
f6c42823
f6d42a23
f6e42c23
f6f42e23
fbc40713
f6040793
00070593
00078513
d1dff0ef
00100793
fef42623
00b00793
fef42423
0b80006f
fe842703
00600793
00f71463
fe042623
fe842783
ff078793
008787b3
fcc7c783
02079e63
fec42783
00078e63
fac42783
00178713
fae42623
02000713
00e78023
0480006f
fac42783
00178713
fae42623
03000713
00e78023
0300006f
fe042623
fe842783
ff078793
008787b3
fcc7c703
fac42783
00178693
fad42623
03070713
0ff77713
00e78023
fe842703
00600793
00f71c63
fac42783
00178713
fae42623
02e00713
00e78023
fe842783
fff78793
fef42423
fe842783
f407d4e3
fac42783
00178713
fae42623
00078023
00000013
09c12083
09812403
09412483
0a010113
00008067
f8010113
06112e23
06812c23
06912a23
08010413
00002497
c9848493
fc040793
00078513
d98fe0ef
fc042883
fc442803
fc842503
fcc42583
fd042603
fd442683
fd842703
fdc42783
0114a023
0104a223
00a4a423
00b4a623
00c4a823
00d4aa23
00e4ac23
00f4ae23
00002797
c4478793
00a00713
00e7a023
00002497
c7448493
fc040793
00078513
d34fe0ef
fc042883
fc442803
fc842503
fcc42583
fd042603
fd442683
fd842703
fdc42783
0114a023
0104a223
00a4a423
00b4a623
00c4a823
00d4aa23
00e4ac23
00f4ae23
00002797
c2078793
00100713
00e7a023
fe042623
1600006f
fec42703
00300793
04f71a63
00002797
bdc78793
00002717
bf470713
00072303
00472883
00872803
00c72503
01072583
01472603
01872683
01c72703
0067a023
0117a223
0107a423
00a7a623
00b7a823
00c7aa23
00d7ac23
00e7ae23
00002497
bac48493
fc040313
00002797
ba078793
0007a883
0047a803
0087a503
00c7a583
0107a603
0147a683
0187a703
01c7a783
fb142023
fb042223
faa42423
fab42623
fac42823
fad42a23
fae42c23
faf42e23
00002797
b1878793
0007a883
0047a803
0087a503
00c7a583
0107a603
0147a683
0187a703
01c7a783
f9142023
f9042223
f8a42423
f8b42623
f8c42823
f8d42a23
f8e42c23
f8f42e23
f8040713
fa040793
00070613
00078593
00030513
f5cfe0ef
fc042883
fc442803
fc842503
fcc42583
fd042603
fd442683
fd842703
fdc42783
0114a023
0104a223
00a4a423
00b4a623
00c4a823
00d4aa23
00e4ac23
00f4ae23
fec42783
00178793
fef42623
fec42703
00500793
e8e7dee3
00002497
ac048493
f8040313
00002797
a9478793
0007a883
0047a803
0087a503
00c7a583
0107a603
0147a683
0187a703
01c7a783
fb142023
fb042223
faa42423
fab42623
fac42823
fad42a23
fae42c23
faf42e23
00002797
a4c78793
0007a883
0047a803
0087a503
00c7a583
0107a603
0147a683
0187a703
01c7a783
fd142023
fd042223
fca42423
fcb42623
fcc42823
fcd42a23
fce42c23
fcf42e23
fc040713
fa040793
00070613
00078593
00030513
e50fe0ef
f8042883
f8442803
f8842503
f8c42583
f9042603
f9442683
f9842703
f9c42783
0114a023
0104a223
00a4a423
00b4a623
00c4a823
00d4aa23
00e4ac23
00f4ae23
00002797
9ec78793
0007a023
00002497
9e048493
f8040793
00078513
a60fe0ef
f8042883
f8442803
f8842503
f8c42583
f9042603
f9442683
f9842703
f9c42783
0714a223
0704a423
06a4a623
06b4a823
06c4aa23
06d4ac23
06e4ae23
08f4a023
00002797
98c78793
00002717
98470713
06472303
06872883
06c72803
07072503
07472583
07872603
07c72683
08072703
0467a223
0517a423
0507a623
04a7a823
04b7aa23
04c7ac23
04d7ae23
06e7a023
00002797
93c78793
00002717
93470713
04472303
04872883
04c72803
05072503
05472583
05872603
05c72683
06072703
0267a223
0317a423
0307a623
02a7a823
02b7aa23
02c7ac23
02d7ae23
04e7a023
00002797
8ec78793
00002717
8e470713
02472303
02872883
02c72803
03072503
03472583
03872603
03c72683
04072703
0067a223
0117a423
0107a623
00a7a823
00b7aa23
00c7ac23
00d7ae23
02e7a023
00002797
89c78793
0807a223
00002797
89078793
0807a423
00002797
88478793
02000713
08e78623
00000013
07c12083
07812403
07412483
08010113
00008067
e5010113
1a112623
1a812423
1a912223
1b010413
00050793
eaf40fa3
fe042423
ee440793
00078513
8c4fe0ef
ebf44703
02f00793
7ae7f063
ebf44703
03900793
78e7ea63
00002797
81878793
ebf44703
08e78623
00002797
80878793
0887a783
16078063
00001797
7f878793
0807a423
00001797
7ec78793
00001717
7e470713
04472303
04872883
04c72803
05072503
05472583
05872603
05c72683
06072703
0667a223
0717a423
0707a623
06a7a823
06b7aa23
06c7ac23
06d7ae23
08e7a023
00001797
79c78793
00001717
79470713
02472303
02872883
02c72803
03072503
03472583
03872603
03c72683
04072703
0467a223
0517a423
0507a623
04a7a823
04b7aa23
04c7ac23
04d7ae23
06e7a023
00001797
74c78793
00001717
74470713
00472303
00872883
00c72803
01072503
01472583
01872603
01c72683
02072703
0267a223
0317a423
0307a623
02a7a823
02b7aa23
02c7ac23
02d7ae23
04e7a023
00001497
6fc48493
e9040793
00078513
f7dfd0ef
e9042883
e9442803
e9842503
e9c42583
ea042603
ea442683
ea842703
eac42783
0114a223
0104a423
00a4a623
00b4a823
00c4aa23
00d4ac23
00e4ae23
02f4a023
00001797
6a878793
0007a023
ebf44783
fd078793
fef42223
00001797
69078793
0007a783
28079a63
00001497
68048493
e9040313
00001797
67478793
0047a883
0087a803
00c7a503
0107a583
0147a603
0187a683
01c7a703
0207a783
e7142823
e7042a23
e6a42c23
e6b42e23
e8c42023
e8d42223
e8e42423
e8f42623
00001797
5ac78793
0007a883
0047a803
0087a503
00c7a583
0107a603
0147a683
0187a703
01c7a783
e5142823
e5042a23
e4a42c23
e4b42e23
e6c42023
e6d42223
e6e42423
e6f42623
e5040713
e7040793
00070613
00078593
00030513
9f0fe0ef
e9042883
e9442803
e9842503
e9c42583
ea042603
ea442683
ea842703
eac42783
0114a223
0104a423
00a4a623
00b4a823
00c4aa23
00d4ac23
00e4ae23
02f4a023
fe442783
eef42223
f0440313
ee442883
ee842803
eec42503
ef042583
ef442603
ef842683
efc42703
f0042783
e5142823
e5042a23
e4a42c23
e4b42e23
e6c42023
e6d42223
e6e42423
e6f42623
00001797
50078793
0007a883
0047a803
0087a503
00c7a583
0107a603
0147a683
0187a703
01c7a783
e7142823
e7042a23
e6a42c23
e6b42e23
e8c42023
e8d42223
e8e42423
e8f42623
e7040713
e5040793
00070613
00078593
00030513
904fe0ef
00001497
4e048493
e5040313
00001797
4d478793
0047a883
0087a803
00c7a503
0107a583
0147a603
0187a683
01c7a703
0207a783
e7142823
e7042a23
e6a42c23
e6b42e23
e8c42023
e8d42223
e8e42423
e8f42623
f0442883
f0842803
f0c42503
f1042583
f1442603
f1842683
f1c42703
f2042783
e9142823
e9042a23
e8a42c23
e8b42e23
eac42023
ead42223
eae42423
eaf42623
e9040713
e7040793
00070613
00078593
00030513
d61fd0ef
e5042883
e5442803
e5842503
e5c42583
e6042603
e6442683
e6842703
e6c42783
0114a223
0104a423
00a4a623
00b4a823
00c4aa23
00d4ac23
00e4ae23
02f4a023
5300006f
00001797
3f078793
0007a703
00700793
50f70e63
00001797
39c78793
0007a883
0047a803
0087a503
00c7a583
0107a603
0147a683
0187a703
01c7a783
ef142223
ef042423
eea42623
eeb42823
eec42a23
eed42c23
eee42e23
f0f42023
fe042623
0f80006f
e5040313
ee442883
ee842803
eec42503
ef042583
ef442603
ef842683
efc42703
f0042783
e7142823
e7042a23
e6a42c23
e6b42e23
e8c42023
e8d42223
e8e42423
e8f42623
00001797
2c878793
0007a883
0047a803
0087a503
00c7a583
0107a603
0147a683
0187a703
01c7a783
e9142823
e9042a23
e8a42c23
e8b42e23
eac42023
ead42223
eae42423
eaf42623
ec440693
e9040713
e7040793
00070613
00078593
00030513
b48fe0ef
e5042883
e5442803
e5842503
e5c42583
e6042603
e6442683
e6842703
e6c42783
ef142223
ef042423
eea42623
eeb42823
eec42a23
eed42c23
eee42e23
f0f42023
fec42783
00178793
fef42623
00001797
29878793
0007a783
fec42703
eef74ee3
e5040793
00078513
b0dfd0ef
e5042883
e5442803
e5842503
e5c42583
e6042603
e6442683
e6842703
e6c42783
ed142223
ed042423
eca42623
ecb42823
ecc42a23
ecd42c23
ece42e23
eef42023
fe442783
ecf42223
f2440313
ee442883
ee842803
eec42503
ef042583
ef442603
ef842683
efc42703
f0042783
e5142823
e5042a23
e4a42c23
e4b42e23
e6c42023
e6d42223
e6e42423
e6f42623
ec442883
ec842803
ecc42503
ed042583
ed442603
ed842683
edc42703
ee042783
e7142823
e7042a23
e6a42c23
e6b42e23
e8c42023
e8d42223
e8e42423
e8f42623
e7040713
e5040793
00070613
00078593
00030513
db9fd0ef
00001497
19448493
e5040313
00001797
18878793
0047a883
0087a803
00c7a503
0107a583
0147a603
0187a683
01c7a703
0207a783
e7142823
e7042a23
e6a42c23
e6b42e23
e8c42023
e8d42223
e8e42423
e8f42623
f2442883
f2842803
f2c42503
f3042583
f3442603
f3842683
f3c42703
f4042783
e9142823
e9042a23
e8a42c23
e8b42e23
eac42023
ead42223
eae42423
eaf42623
e9040713
e7040793
00070613
00078593
00030513
a15fd0ef
e5042883
e5442803
e5842503
e5c42583
e6042603
e6442683
e6842703
e6c42783
0114a223
0104a423
00a4a623
00b4a823
00c4aa23
00d4ac23
00e4ae23
02f4a023
00001797
0a878793
0007a783
00178713
00001797
09878793
00e7a023
1c80006f
ebf44703
02e00793
02f71c63
00001797
07c78793
0007a783
1a079863
00001797
06c78793
00100713
00e7a023
00001797
05c78793
02e00713
08e78623
18c0006f
ebf44703
00d00793
16f71463
00001797
03c78793
03b00713
08e78623
00001797
02c78793
00001717
02470713
04472303
04872883
04c72803
05072503
05472583
05872603
05c72683
06072703
0667a223
0717a423
0707a623
06a7a823
06b7aa23
06c7ac23
06d7ae23
08e7a023
00001797
fdc78793
00001717
fd470713
02472303
02872883
02c72803
03072503
03472583
03872603
03c72683
04072703
0467a223
0517a423
0507a623
04a7a823
04b7aa23
04c7ac23
04d7ae23
06e7a023
00001797
f8c78793
00001717
f8470713
00472303
00872883
00c72803
01072503
01472583
01872603
01c72683
02072703
0267a223
0317a423
0307a623
02a7a823
02b7aa23
02c7ac23
02d7ae23
04e7a023
00001497
f3c48493
e5040793
00078513
fbcfd0ef
e5042883
e5442803
e5842503
e5c42583
e6042603
e6442683
e6842703
e6c42783
0114a223
0104a423
00a4a623
00b4a823
00c4aa23
00d4ac23
00e4ae23
02f4a023
00001797
ee878793
0007a023
01c0006f
ebf44703
07200793
00f71863
9a0ff0ef
0080006f
00000013
ebf44703
02b00793
02f70463
ebf44703
02d00793
00f70e63
ebf44703
02a00793
00f70863
ebf44703
02f00793
60f71a63
00001797
e9078793
ebf44703
08e78623
ebf44703
02b00793
0ef71c63
00001497
e7448493
e5040313
00001797
e6878793
0047a883
0087a803
00c7a503
0107a583
0147a603
0187a683
01c7a703
0207a783
e7142823
e7042a23
e6a42c23
e6b42e23
e8c42023
e8d42223
e8e42423
e8f42623
00001797
e2078793
0247a883
0287a803
02c7a503
0307a583
0347a603
0387a683
03c7a703
0407a783
e9142823
e9042a23
e8a42c23
e8b42e23
eac42023
ead42223
eae42423
eaf42623
e9040713
e7040793
00070613
00078593
00030513
eecfd0ef
e5042883
e5442803
e5842503
e5c42583
e6042603
e6442683
e6842703
e6c42783
0114a223
0104a423
00a4a623
00b4a823
00c4aa23
00d4ac23
00e4ae23
02f4a023
ebf44703
02d00793
0ef71c63
00001497
d7448493
e5040313
00001797
d6878793
0247a883
0287a803
02c7a503
0307a583
0347a603
0387a683
03c7a703
0407a783
e7142823
e7042a23
e6a42c23
e6b42e23
e8c42023
e8d42223
e8e42423
e8f42623
00001797
d2078793
0047a883
0087a803
00c7a503
0107a583
0147a603
0187a683
01c7a703
0207a783
e9142823
e9042a23
e8a42c23
e8b42e23
eac42023
ead42223
eae42423
eaf42623
e9040713
e7040793
00070613
00078593
00030513
f68fd0ef
e5042883
e5442803
e5842503
e5c42583
e6042603
e6442683
e6842703
e6c42783
0114a223
0104a423
00a4a623
00b4a823
00c4aa23
00d4ac23
00e4ae23
02f4a023
ebf44703
02a00793
1af71063
f4440313
00001797
c7078793
0047a883
0087a803
00c7a503
0107a583
0147a603
0187a683
01c7a703
0207a783
e5142823
e5042a23
e4a42c23
e4b42e23
e6c42023
e6d42223
e6e42423
e6f42623
00001797
c2878793
0247a883
0287a803
02c7a503
0307a583
0347a603
0387a683
03c7a703
0407a783
e7142823
e7042a23
e6a42c23
e6b42e23
e8c42023
e8d42223
e8e42423
e8f42623
e7040713
e5040793
00070613
00078593
00030513
fecfd0ef
00001497
bc848493
e5040313
f4442883
f4842803
f4c42503
f5042583
f5442603
f5842683
f5c42703
f6042783
e7142823
e7042a23
e6a42c23
e6b42e23
e8c42023
e8d42223
e8e42423
e8f42623
00001797
b3c78793
0007a883
0047a803
0087a503
00c7a583
0107a603
0147a683
0187a703
01c7a783
e9142823
e9042a23
e8a42c23
e8b42e23
eac42023
ead42223
eae42423
eaf42623
ee440693
e9040713
e7040793
00070613
00078593
00030513
b7dfd0ef
e5042883
e5442803
e5842503
e5c42583
e6042603
e6442683
e6842703
e6c42783
0114a223
0104a423
00a4a623
00b4a823
00c4aa23
00d4ac23
00e4ae23
02f4a023
ebf44703
02f00793
1af71063
f6440313
00001797
ac878793
0247a883
0287a803
02c7a503
0307a583
0347a603
0387a683
03c7a703
0407a783
e5142823
e5042a23
e4a42c23
e4b42e23
e6c42023
e6d42223
e6e42423
e6f42623
00001797
a4078793
0007a883
0047a803
0087a503
00c7a583
0107a603
0147a683
0187a703
01c7a783
e7142823
e7042a23
e6a42c23
e6b42e23
e8c42023
e8d42223
e8e42423
e8f42623
e7040713
e5040793
00070613
00078593
00030513
e44fd0ef
00001497
a2048493
e5040313
f6442883
f6842803
f6c42503
f7042583
f7442603
f7842683
f7c42703
f8042783
e7142823
e7042a23
e6a42c23
e6b42e23
e8c42023
e8d42223
e8e42423
e8f42623
00001797
9d478793
0047a883
0087a803
00c7a503
0107a583
0147a603
0187a683
01c7a703
0207a783
e9142823
e9042a23
e8a42c23
e8b42e23
eac42023
ead42223
eae42423
eaf42623
ee440693
e9040713
e7040793
00070613
00078593
00030513
9d5fd0ef
e5042883
e5442803
e5842503
e5c42583
e6042603
e6442683
e6842703
e6c42783
0114a223
0104a423
00a4a623
00b4a823
00c4aa23
00d4ac23
00e4ae23
02f4a023
00001797
93078793
00001717
92870713
04472303
04872883
04c72803
05072503
05472583
05872603
05c72683
06072703
0267a223
0317a423
0307a623
02a7a823
02b7aa23
02c7ac23
02d7ae23
04e7a023
00001797
8e078793
00001717
8d870713
06472303
06872883
06c72803
07072503
07472583
07872603
07c72683
08072703
0467a223
0517a423
0507a623
04a7a823
04b7aa23
04c7ac23
04d7ae23
06e7a023
00001797
89078793
00100713
08e7a423
ebf44703
07300793
14f71e63
f8440313
00001797
87078793
0047a883
0087a803
00c7a503
0107a583
0147a603
0187a683
01c7a703
0207a783
e5142823
e5042a23
e4a42c23
e4b42e23
e6c42023
e6d42223
e6e42423
e6f42623
00000797
7e878793
0007a883
0047a803
0087a503
00c7a583
0107a603
0147a683
0187a703
01c7a783
e7142823
e7042a23
e6a42c23
e6b42e23
e8c42023
e8d42223
e8e42423
e8f42623
e7040713
e5040793
00070613
00078593
00030513
becfd0ef
00000497
7c848493
e5040313
f8442883
f8842803
f8c42503
f9042583
f9442603
f9842683
f9c42703
fa042783
e7142823
e7042a23
e6a42c23
e6b42e23
e8c42023
e8d42223
e8e42423
e8f42623
e7040793
00078593
00030513
864fe0ef
e5042883
e5442803
e5842503
e5c42583
e6042603
e6442683
e6842703
e6c42783
0114a223
0104a423
00a4a623
00b4a823
00c4aa23
00d4ac23
00e4ae23
02f4a023
00000797
72c78793
00100713
08e7a423
00000797
71c78793
0847a783
02078463
ebf44703
00d00793
00f70e63
ebf44703
00a00793
00f70863
00000797
6f478793
0807a223
00000797
6e878793
0047a883
0087a803
00c7a503
0107a583
0147a603
0187a683
01c7a703
0207a783
ef142223
ef042423
eea42623
eeb42823
eec42a23
eed42c23
eee42e23
f0f42023
ee442883
ee842803
eec42503
ef042583
ef442603
ef842683
efc42703
f0042783
e5142823
e5042a23
e4a42c23
e4b42e23
e6c42023
e6d42223
e6e42423
e6f42623
e5040793
00078513
cd4fd0ef
00050793
0e078663
fa440793
00078513
ed5fc0ef
e5040313
fa442883
fa842803
fac42503
fb042583
fb442603
fb842683
fbc42703
fc042783
e7142823
e7042a23
e6a42c23
e6b42e23
e8c42023
e8d42223
e8e42423
e8f42623
ee442883
ee842803
eec42503
ef042583
ef442603
ef842683
efc42703
f0042783
e9142823
e9042a23
e8a42c23
e8b42e23
eac42023
ead42223
eae42423
eaf42623
e9040713
e7040793
00070613
00078593
00030513
84cfd0ef
e5042883
e5442803
e5842503
e5c42583
e6042603
e6442683
e6842703
e6c42783
ef142223
ef042423
eea42623
eeb42823
eec42a23
eed42c23
eee42e23
f0f42023
fc440313
ee442883
ee842803
eec42503
ef042583
ef442603
ef842683
efc42703
f0042783
e5142823
e5042a23
e4a42c23
e4b42e23
e6c42023
e6d42223
e6e42423
e6f42623
00000797
50078793
0007a883
0047a803
0087a503
00c7a583
0107a603
0147a683
0187a703
01c7a783
e7142823
e7042a23
e6a42c23
e6b42e23
e8c42023
e8d42223
e8e42423
e8f42623
e7040713
e5040793
00070613
00078593
00030513
f69fc0ef
fc442883
fc842803
fcc42503
fd042583
fd442603
fd842683
fdc42703
fe042783
e5142823
e5042a23
e4a42c23
e4b42e23
e6c42023
e6d42223
e6e42423
e6f42623
e5040793
00078513
af4fd0ef
00050793
06079463
00000797
46c78793
00100713
08e7a223
00000497
45c48493
e5040793
00078513
cddfc0ef
e5042883
e5442803
e5842503
e5c42583
e6042603
e6442683
e6842703
e6c42783
0114a223
0104a423
00a4a623
00b4a823
00c4aa23
00d4ac23
00e4ae23
02f4a023
00000013
1ac12083
1a812403
1a412483
1b010113
00008067
f8010113
06112e23
06812c23
08010413
00000797
35c78793
0007a023
ea8fe0ef
00000517
29850513
bd0fe0ef
00000797
3c478793
0647a883
0687a803
06c7a503
0707a583
0747a603
0787a683
07c7a703
0807a783
f9142023
f9042223
f8a42423
f8b42623
f8c42823
f8d42a23
f8e42c23
f8f42e23
fa040713
f8040793
00070593
00078513
bb4fe0ef
00000797
36878793
0447a883
0487a803
04c7a503
0507a583
0547a603
0587a683
05c7a703
0607a783
f9142023
f9042223
f8a42423
f8b42623
f8c42823
f8d42a23
f8e42c23
f8f42e23
fa040793
01478713
f8040793
00070593
00078513
b54fe0ef
00000797
30878793
0247a883
0287a803
02c7a503
0307a583
0347a603
0387a683
03c7a703
0407a783
f9142023
f9042223
f8a42423
f8b42623
f8c42823
f8d42a23
f8e42c23
f8f42e23
fa040793
02878713
f8040793
00070593
00078513
af4fe0ef
00000797
2a878793
0047a883
0087a803
00c7a503
0107a583
0147a603
0187a683
01c7a703
0207a783
f9142023
f9042223
f8a42423
f8b42623
f8c42823
f8d42a23
f8e42c23
f8f42e23
fa040793
03c78713
f8040793
00070593
00078513
a94fe0ef
00000517
13050513
a48fe0ef
00000517
13c50513
a3cfe0ef
00000517
16450513
a30fe0ef
fa040793
00078513
a24fe0ef
00000517
15450513
a18fe0ef
00000517
14c50513
a0cfe0ef
fa040793
01478793
00078513
9fcfe0ef
00000517
12c50513
9f0fe0ef
00000517
12c50513
9e4fe0ef
fa040793
02878793
00078513
9d4fe0ef
00000517
10450513
9c8fe0ef
00000517
10c50513
9bcfe0ef
fa040793
03c78793
00078513
9acfe0ef
00000517
0dc50513
9a0fe0ef
00000797
19478793
0847a783
00078863
00000517
0dc50513
984fe0ef
00000517
0b450513
978fe0ef
00000517
0d850513
96cfe0ef
00100593
00000517
1e850513
825fc0ef
8f5fc0ef
00050793
00078513
8e9fe0ef
d7dff06f
ffff0000
2d524159
636c6143
74616c75
5320726f
74726174
20676e69
2e2e7075
000a0d2e
3d3d3d3d
3d3d3d3d
3d3d3d3d
3d3d3d3d
3d3d3d3d
00000000
2d524159
636f7250
6f737365
70412072
63696c70
6f697461
6544206e
203a6f6d
204e5052
636c6143
74616c75
0d0a726f
00000000
203a5409
00000000
00000d0a
203a5a09
00000000
203a5909
00000000
203a5809
00000000
4e524157
3a474e49
65764f20
6f6c6672
00000077
7473614c
79654b20
0000203a
80000000
