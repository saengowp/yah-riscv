800000b7
00000137
10010113
00010183
fe018ae3
0000c203
00f27213
001202b3
02028293
00328023
00120213
00f27213
00408023
0000c283
0f02f293
0042d293
fe521ae3
00110113
fc5ff06f
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
6c6c6548
6f57206f
0d646c72
0000000a
