00007137
00007437
0040006f
fe010113
00112e23
00812c23
02010413
15c00793
fef42623
fec42503
0e4000ef
00050793
00078593
fec42503
018000ef
00000013
01c12083
01812403
02010113
00008067
fd010113
02812623
03010413
fca42e23
fcb42c23
08c0006f
16c02783
0007c783
fef407a3
fef44783
0047d793
fef40723
fef44783
00f7f793
fef406a3
fed44783
00178793
0ff7f793
00f7f793
fef40623
fec44703
fee44783
00f71463
0440006f
16c02703
fed44783
02078793
00f707b3
fdc42703
00074703
00e78023
16c02783
fec44703
00e78023
fdc42783
00178793
fcf42e23
fd842783
fff78793
fcf42c23
fd842783
f6079ae3
00000013
00000013
02c12403
03010113
00008067
fd010113
02812623
03010413
fca42e23
fe042623
01c0006f
fec42783
00178793
fef42623
fdc42783
00178793
fcf42e23
fdc42783
0007c783
fe0790e3
fec42783
00078513
02c12403
03010113
00008067
6c6c6548
6f57206f
21646c72
00000000
80000000
