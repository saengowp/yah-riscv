00007137
00007437
00000517
1a850513
00050067
fd010113
02812623
03010413
fca42e23
fcb42c23
0980006f
21000793
0007a783
0007c783
fef407a3
fef44783
0047d793
fef40723
fef44783
00f7f793
fef406a3
fed44783
00178793
0ff7f793
00f7f793
fef40623
fec44703
fee44783
00f71463
04c0006f
21000793
0007a703
fed44783
02078793
00f707b3
fdc42703
00074703
00e78023
21000793
0007a783
fec44703
00e78023
fdc42783
00178793
fcf42e23
fd842783
fff78793
fcf42c23
fd842783
f60794e3
00000013
00000013
02c12403
03010113
00008067
fe010113
00812e23
02010413
21000793
0007a783
0017c783
fef407a3
fef44783
00f7f793
fef407a3
fef44703
21400793
0007a783
fcf70ce3
21000793
0007a703
21400793
0007a783
01078793
00f707b3
0007c783
fef40723
21400793
0007a783
00178793
00f7f713
21400793
00e7a023
fee44783
00078513
01c12403
02010113
00008067
fd010113
02812623
03010413
fca42e23
fe042623
01c0006f
fec42783
00178793
fef42623
fdc42783
00178793
fcf42e23
fdc42783
0007c783
fe0790e3
fec42783
00078513
02c12403
03010113
00008067
fe010113
00112e23
00812c23
02010413
20000793
fef42623
fec42503
f95ff0ef
00050793
00078593
fec42503
e39ff0ef
efdff0ef
00050793
fef405a3
feb40793
00100593
00078513
e1dff0ef
fe5ff06f
6c6c6548
6f57206f
21646c72
00000a0d
80000000
