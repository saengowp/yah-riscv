2a000113
20400513
0a4000ef
000024b7
00000913
02000993
0c8000ef
00050a13
0fc000ef
02000513
ff4508e3
00d00513
ff4504e3
00a00513
ff4500e3
00a00593
fd0a0513
00a5e463
0180006f
00500593
f9fa0513
02a5ea63
00a50513
0040006f
00491913
00a96933
ffc98993
fa0996e3
0124a023
00448493
02000993
24e00513
02c000ef
f95ff06f
04a00513
01451a63
26400513
018000ef
00002537
00050067
28800513
008000ef
f71ff06f
00112023
00912223
00810113
00050493
00048503
00050863
058000ef
00148493
ff1ff06f
ff810113
00012083
00412483
00008067
00112023
00410113
074000ef
20000e13
000e2383
fe750ae3
01068313
00730333
00034503
00138393
00f3f393
007e2023
ffc10113
00012083
00008067
00112023
00a12223
00810113
034000ef
ffc10113
00012503
02068293
00c282b3
00a28023
00160313
00668023
014000ef
fec59ee3
ffc10113
00012083
00008067
800006b7
0006a283
00028513
00028593
00028613
00855513
0045d593
00f57513
00f5f593
00f67613
00008067
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
2d484159
43534952
6f432056
42206572
6c746f6f
6564616f
4c0a0d72
65747369
676e696e
206f7420
676f7270
206d6172
0d786568
6174530a
6e697472
74612067
32783020
0d303030
0a0d000a
64726f57
6b636120
6c776f6e
65676465
000a0d64
204a0a0d
65636552
64657669
6f43202e
6f72746e
7254206c
66736e61
2e2e7265
000a0d2e
61766e49
2064696c
72616863
63657220
65766965
000a0d64
00000000
